/* target_ipi.cdl */

import("tIPI.cdl");

