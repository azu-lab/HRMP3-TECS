/*
 *		C言語で記述されたアプリケーションから，TECSベースの実行時間分布
 *		集計サービスを呼び出すためのアダプタ用セルタイプの定義
 * 
 *  $Id: tHistogramAdapter.cdl 3234 2021-10-24 13:13:34Z ertl-hiro $
 */
[singleton, active]
celltype tHistogramAdapter {
	call	sHistogram		cHistogram[];
};
