/*
 *		C言語で記述されたアプリケーションから，TECSベースのテストプログ
 *		ラム用サービスを呼び出すためのアダプタ用セルタイプの定義
 *
 *  $Id: tTestServiceAdapter.cdl 3234 2021-10-24 13:13:34Z ertl-hiro $
 */
[singleton, active]
celltype tTestServiceAdapter {
	call	sTestService	cTestService;
};
