/*
 *  TOPPERS Software
 *      Toyohashi Open Platform for Embedded Real-Time Systems
 * 
 *  Copyright (C) 2015 by Ushio Laboratory
 *              Graduate School of Engineering Science, Osaka Univ., JAPAN
 *  Copyright (C) 2015,2016 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 * 
 *  上記著作権者は，以下の(1)〜(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 * 
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 * 
 *  $Id: tSysLog.cdl 3234 2021-10-24 13:13:34Z ertl-hiro $
 */

/*
 *		システムログ機能のコンポーネント記述ファイル
 */

/*
 *  システムログ機能に関する定義
 */
import_C("syssvc/syslog.h");

/*
 *  低レベル出力のシグニチャ
 */
signature sPutLog {
	void	putChar([in] char c);
};

/*
 *  システムログ機能のシグニチャ
 */
signature sSysLog {
	/*
	 *  ログ情報の出力
	 */
	ER		write([in] uint_t priority, [in] const SYSLOG *p_syslog);

	/*
	 *  ログバッファからのログ情報の読出し
	 */
	ER_UINT	read([out] SYSLOG *p_syslog);

	/*
	 *  出力すべきログ情報の重要度の設定
	 */
	ER		mask([in] uint_t logMask, [in] uint_t lowMask);

	/*
	 *  ログバッファの状態参照
	 */
	ER		refer([out] T_SYSLOG_RLOG *pk_rlog);

	/*
	 *  低レベル出力によるすべてのログ情報の出力
	 */
	ER		flush(void);
};

/*
 *  システムログ機能のセルタイプ
 */
[singleton]
celltype tSysLog {
	entry	sSysLog		eSysLog;
	call	sPutLog		cPutLog;		/* 低レベル出力との接続 */

	attr {
		uint_t	logBufferSize;			/* ログバッファサイズ */
		uint_t	initLogMask = C_EXP("LOG_UPTO(LOG_DEBUG)");
										/* ログバッファに記録すべき重要度 */
		uint_t	initLowMask = C_EXP("LOG_UPTO(LOG_EMERG)");
									   	/* 低レベル出力すべき重要度 */
	};
	var {
		[size_is(logBufferSize)] SYSLOG	*logBuffer;	/* ログバッファ */
		uint_t	count = 0;				/* ログバッファ中のログの数 */
		uint_t	head = 0;				/* 先頭のログの格納位置 */
		uint_t	tail = 0;				/* 次のログの格納位置 */
		uint_t	lost = 0;				/* 失われたログの数 */
		uint_t	logMask = initLogMask;	/* ログバッファに記録すべき重要度 */
		uint_t	lowMask = initLowMask;	/* 低レベル出力すべき重要度 */
	};
};
