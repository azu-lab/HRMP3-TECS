import(<kernel.cdl>);

region rKernelDomain{
region rProcessor1Migratable{
    cell tTask Task1 {
        /* 呼び口の結合 */
        cTaskBody = rProcessor1Migratable::Exc08.eSampleTask[0];
        /* 属性の設定 */
        priority = C_EXP("MID_PRIORITY");
        stackSize = C_EXP("STACK_SIZE");
    };
    
    cell tTask Task2 {
        /* 呼び口の結合 */
        cTaskBody = rProcessor1Migratable::Exc08.eSampleTask[1];
        /* 属性の設定 */
        priority = C_EXP("MID_PRIORITY");
        stackSize = C_EXP("STACK_SIZE");
    };
};

[domain(HRMP, "user")]
region rUserDomain1{
	[class(HRMP,"CLS_PRC1")]
	region rProcessor1Only{
		cell tSample Sample1{
			cSample = Sample2.eSample;
		};

		cell tSample Sample1{
			cSample = Sample2.eSample;
		};
	};
	[class(HRMP, "CLS_PRC2")]
	region rProcessor2Only{
		cell tSample Sample2{
			cSample = Sample2.eSample;
		};
	};
	[class(HRMP, "CLS_PRC3")]
	region rProcessor3Only{
		cell tSample Sample2{
			cSample = Sample2.eSample;
		};
	};	
};

[domain(HRMP,"user")]
region rUserDomain2{
	[class(HRMP, "CLS_ALL_PRC1")]
	region rProcessor1Mig{
		cell tSample Sample3{
			cSample = Sample2.eSample;
		};
	};	
};
