/* tSIOPortZyboZ7.cdl */ 

// import_C("target_syssvc.h");
import_C("zybo_z7.h");
import_C("zynq7000.h");

import("tXUartPs.cdl");

celltype tSIOPortZyboZ7Main{
	/*
	 *  シリアルインタフェースドライバとの結合
	 */
	[inline] entry		sSIOPort	eSIOPort;
	[optional] call		siSIOCBR	ciSIOCBR;

	/*
	 *  SIOドライバとの結合
	 */
	call			sSIOPort	cSIOPort;
	[inline] entry	siSIOCBR	eiSIOCBR;

	/*
	 *  割込み要求ライン操作のための結合
	 */
	call	sInterruptRequest	cInterruptRequest;
};

/*
 *  シリアルインタフェースドライバのターゲット依存部（複合コンポーネン
 *  ト）のセルタイプ
 */
[active]
composite tSIOPortZyboZ7 {
	/*
	 *  シリアルインタフェースドライバとの結合
	 */
	entry				sSIOPort	eSIOPort;
	[optional] call		siSIOCBR	ciSIOCBR;

	/*
	 *  属性の定義
	 */
	attr {
		uintptr_t	baseAddress;														/* ベースアドレス */
		INTNO		interruptNumber;													/* 割込み番号 */
		PRI			isrPriority = C_EXP("1");				/* ISR優先度 */
		PRI			interruptPriority = C_EXP("(-4)");	/* 割込み優先度 */
		/*
		PRI			isrPriority = C_EXP("ISRPRI_SIO");				/* ISR優先度 *
		PRI			interruptPriority = C_EXP("INTPRI_SIO");	/* 割込み優先度 *
		*/

		uint16_t		baudgen = C_EXP("XUARTPS_BAUDGEN_115K"); // 8bit, non-parity, 1stop-bit
		uint8_t			bauddiv = C_EXP("XUARTPS_BAUDDIV_115K"); // 115K baud
		uint16_t		mode    = C_EXP("XUARTPS_MR_CHARLEN_8 | XUARTPS_MR_PARITY_NONE | XUARTPS_MR_STOPBIT_1");    // 115K baud
		/*
		uint16_t		baudgen = C_EXP("SIO_XUARTPS_BAUDGEN"); // 8bit, non-parity, 1stop-bit
		uint8_t			bauddiv = C_EXP("SIO_XUARTPS_BAUDDIV"); // 115K baud
		uint16_t		mode    = C_EXP("SIO_XUARTPS_MODE");    // 115K baud
		*/
	};

	/*
	 *  SIOドライバ
	 */
	cell tXUartPs XUartPs {
		baseAddress = composite.baseAddress;
		baudgen     = composite.baudgen;
		bauddiv     = composite.bauddiv;
		mode        = composite.mode;
		ciSIOCBR    = SIOPortMain.eiSIOCBR;
	};
	
	/*
	 *  シリアルインタフェースドライバのターゲット依存部の本体
	 */
	cell tSIOPortZyboZ7Main SIOPortMain {
		ciSIOCBR          => composite.ciSIOCBR;
		cSIOPort          = XUartPs.eSIOPort;
		cInterruptRequest = InterruptRequest.eInterruptRequest;
	};
	composite.eSIOPort => SIOPortMain.eSIOPort;

	/*
	 *  SIOの割込みサービスルーチンと割込み要求ライン
	 */
	cell tISR ISRInstance {
		interruptNumber = composite.interruptNumber;
		isrPriority     = composite.isrPriority;
		ciISRBody       = XUartPs.eiISR;
	};
	cell tInterruptRequest InterruptRequest {
		interruptNumber   = composite.interruptNumber;
		interruptPriority = composite.interruptPriority;
	};

  /*
   * 終了処理ルーチン
   */
  cell tTerminateRoutine Terminate {
      cTerminateRoutineBody = XUartPs.eTerminate;
  };
};

// region rOutOfDomain{
region rKernelDomain {
// region rProcessor1Migratable {
region rProcessor1Only {

    /*
     *  シリアルインタフェースドライバのターゲット依存部のプロトタイプ
     */
    [prototype]
        cell tSIOPortZyboZ7 SIOPortTarget1 {
        /* 属性の設定 */
        baseAddress     = C_EXP("ZYNQ_UART1_BASE");
        interruptNumber = C_EXP("ZYNQ_UART1_IRQ");
        /*
        baseAddress     = C_EXP("SIO_XUARTPS_BASE");
        interruptNumber = C_EXP("INTNO_SIO");
        */
    	};
    };

};