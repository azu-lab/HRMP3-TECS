/*
 *      サンプルプログラム(2)のコンポーネント記述ファイル
 *
 *  $Id: tTest_sample.cdl 869 2018-01-04 10:44:46Z ertl-hiro $
 */

/*
 *  カーネルオブジェクトの定義
 */
import(<kernel.cdl>);

/*
 *  ターゲット非依存のセルタイプの定義
 */
import("syssvc/tSerialPort.cdl");
import("syssvc/tSerialAdapter.cdl");
import("syssvc/tSysLog.cdl");
import("syssvc/tSysLogAdapter.cdl");
import("syssvc/tLogTask.cdl");
import("syssvc/tBanner.cdl");

/*
 *  ターゲット依存部の取り込み
 */
import("target.cdl");

/*
 *  サンプルプログラムのC言語ヘッダファイルの取り込み
 */
import_C("tTestSample.h");

// RPC の定義をりこむ 
import( "rpc.cdl" );
import( "tDataqueueOWChannel.cdl" );

/*
 *      システムログ機能のアダプタの組上げ記述
 *
 *  システムログ機能のアダプタは，C言語で記述されたコードから，TECSベー
 *  スのシステムログ機能を呼び出すためのセルである．システムログ機能の
 *  サービスコール（syslog，syslog_0〜syslog_5，t_perrorを含む）を呼び
 *  出さない場合には，以下のセルの組上げ記述を削除してよい．
 */
region rKernelDomain{
    region rProcessor1Migratable {
        cell tSysLogAdapter SysLogAdapter {
            cSysLog = rProcessor1Migratable::SysLog.eSysLog;
        };

        /*
        *       シリアルインタフェースドライバのアダプタの組上げ記述
        *
        *  シリアルインタフェースドライバのアダプタは，C言語で記述されたコー
        *  ドから，TECSベースのシリアルインタフェースドライバを呼び出すための
        *  セルである．シリアルインタフェースドライバのサービスコールを呼び出
        *  さない場合には，以下のセルの組上げ記述を削除してよい．
        */
        cell tSerialAdapter SerialAdapter {
            cSerialPort[0] = rProcessor1Migratable::SerialPort1.eSerialPort;
        };
    };
};

/*
 *  これ以降のセルは，カーネルドメイン内に含める
 */
region rKernelDomain {
    region rProcessor1Migratable {

        /*
        *       システムログ機能の組上げ記述
        *
        *  システムログ機能を外す場合には，以下のセルの組上げ記述を削除し，コ
        *  ンパイルオプションに-DTOPPERS_OMIT_SYSLOGを追加すればよい．ただし，
        *  システムログタスクはシステムログ機能を使用するため，それも外すこと
        *  が必要である．また，システムログ機能のアダプタも外さなければならな
        *  い．tecsgenが警告メッセージを出すが，無視してよい．
        */
        cell tSysLog SysLog {
            logBufferSize = 32;                 /* ログバッファのサイズ */
            initLogMask = C_EXP("LOG_UPTO(LOG_NOTICE)");
                                                /* ログバッファに記録すべき重要度 */
            initLowMask = C_EXP("LOG_UPTO(LOG_EMERG)");
                                                /* 低レベル出力すべき重要度 */
            /* 低レベル出力との結合 */
            cPutLog = rProcessor1Only::PutLogTarget.ePutLog;
        };

        /*
        *       シリアルインタフェースドライバの組上げ記述
        *
        *  シリアルインタフェースドライバを外す場合には，以下のセルの組上げ記
        *  述を削除すればよい．ただし，システムログタスクはシリアルインタフェー
        *  スドライバを使用するため，それも外すことが必要である．また，シリア
        *  ルインタフェースドライバのアダプタも外さなければならない．
        */
        cell tSerialPort SerialPort1 {
            receiveBufferSize = 256;            /* 受信バッファのサイズ */
            sendBufferSize    = 256;            /* 送信バッファのサイズ */

            /* ターゲット依存部との結合 */
            // cSIOPort = SIOPortTarget1.eSIOPort;
            // eiSIOCBR <= SIOPortTarget1.ciSIOCBR;    /* コールバック */
            cSIOPort = rKernelDomain::rProcessor1Only::SIOPortTarget1.eSIOPort;
            eiSIOCBR <= rKernelDomain::rProcessor1Only::SIOPortTarget1.ciSIOCBR;    /* コールバック */
        };

        /*
        *       システムログタスクの組上げ記述
        *
        *  システムログタスクを外す場合には，以下のセルの組上げ記述を削除すれ
        *  ばよい．
        */
        cell tLogTask LogTask {
            priority  = 3;                  /* システムログタスクの優先度 */
            stackSize = LogTaskStackSize;   /* システムログタスクのスタックサイズ */

            /* シリアルインタフェースドライバとの結合 */
            cSerialPort        = SerialPort1.eSerialPort;
            cnSerialPortManage = SerialPort1.enSerialPortManage;

            /* システムログ機能との結合 */
            cSysLog = SysLog.eSysLog;

            /* 低レベル出力との結合 */
            cPutLog = rProcessor1Only::PutLogTarget.ePutLog;
        };

        /*
        *       カーネル起動メッセージ出力の組上げ記述
        *
        *  カーネル起動メッセージの出力を外す場合には，以下のセルの組上げ記述
        *  を削除すればよい．
        */
        cell tBanner Banner {
            /* 属性の設定 */
            targetName      = BannerTargetName;
            copyrightNotice = BannerCopyrightNotice;
        };
    };
};

/*
 *      サンプルプログラムのセルタイプの定義
 */
// [singleton]      // HRMP3 版では singleton ではない
celltype tTestSample {
    require tKernel.eKernel;            /* 呼び口名なし（例：delay）*/
    /*require cKernel = tKernel.eKernel;/* 呼び口名あり（例：cKernel_delay）*/
    require ciKernel = tKernel.eiKernel;/* 呼び口名あり（例：ciKernel_）*/

    call sTask          cTask[2];   /* タスク操作 */

    call sSerialPort    cSerialPort;    /* シリアルドライバとの接続 */
    call sSysLog        cSysLog;        /* システムログ機能との接続 */
    
    entry sTaskBody     eMainTask;      /* Mainタスク */
    entry sTaskBody     eMotor1;    /* モータを模したタスク(PRC1) */
    entry sTaskBody     eMotor2;    /* モータを模したタスク(PRC2) */
    // entry sTaskBody     eDataAcqu1;    /* リアルタイム通信を模したタスク(PRC1) */
    // entry sTaskBody     eDataAcqu2;    /* リアルタイム通信を模したタスク(PRC2) */
};

/*
 *      組み上げ記述
 */
[domain(HRMP, "user")]
region rUserDomain1{
    [class(HRMP,"CLS_PRC1")]
    region rProcessor1Only{
        cell tTask DataAcqu1 {
            /* 呼び口の結合 */
            cTaskBody = rUserDomain1::rProcessor2Only::Motor1.eTask;
            /* 属性の設定 */
            priority = C_EXP("MID_PRIORITY");
            stackSize = C_EXP("STACK_SIZE");
        };
    };
    [class(HRMP,"CLS_PRC2")]
    region rProcessor2Only{
        cell tTask Motor1 {
            /* 呼び口の結合 */
            cTaskBody = rKernelDomain::rProcessor1Migratable::TestSample.eMotor1;
            /* 属性の設定 */
            priority = C_EXP("MID_PRIORITY");
            stackSize = C_EXP("STACK_SIZE");
        };
    };        
};

[domain(HRMP, "user")]
region rUserDomain2{
    [class(HRMP,"CLS_PRC1")]
    region rProcessor1Only{
        cell tTask DataAcqu2 {
            /* 呼び口の結合 */
            cTaskBody = rUserDomain2::rProcessor2Only::Motor2.eTask;
            /* 属性の設定 */
            priority = C_EXP("MID_PRIORITY");
            stackSize = C_EXP("STACK_SIZE");
        };
    };
    [class(HRMP,"CLS_PRC2")]
    region rProcessor2Only{
        cell tTask Motor2 {
            /* 呼び口の結合 */
            cTaskBody = rKernelDomain::rProcessor1Migratable::TestSample.eMotor2;
            /* 属性の設定 */
            priority = C_EXP("MID_PRIORITY");
            stackSize = C_EXP("STACK_SIZE");
        };
    };
};

region rKernelDomain{
    region rProcessor1Migratable {
        cell tTask MainTask {
            /* 呼び口の結合 */
            cTaskBody = TestSample.eMainTask;
            /* 属性の設定 */
            attribute = C_EXP("TA_ACT");
            priority = C_EXP("MAIN_PRIORITY");
            stackSize = C_EXP("STACK_SIZE");
        };
    
        cell tTestSample TestSample{
            /* 呼び口の結合 */
            cTask[0] = rUserDomain1::rProcessor1Only::DataAcqu1.eTask;
            cTask[1] = rUserDomain2::rProcessor1Only::DataAcqu2.eTask;

            cSerialPort = rProcessor1Migratable::SerialPort1.eSerialPort;
            cSysLog     = rProcessor1Migratable::SysLog.eSysLog;
        };
    };

    cell tKernel Kernel {
    };
};
